/********************MangoMIPS32*******************
Filename:	CP0.v
Author:		RickyTino
Version:	Unreleased
**************************************************/
`include "Defines.v"

module CP0
(
    input  wire  clk,
    input  wire  rst

);

endmodule